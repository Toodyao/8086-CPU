module ad_control(BHE, A0, in_ad, out_odd, out_even);

input BHE, A0;
input[15:0] in_ad;
output[7:0] out_odd, out_even;

always @(BHE or A0)
begin

end

endmodule
